module Dache(
    input dbus_req_t t_dreq,
    output dbus_resp_t cache_dresp,
);
    
    endmodule
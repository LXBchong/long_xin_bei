`include "common.svh"
`include "instr.svh"

module exhandler(
    
);

endmodule
`include "def.svh"


module Dache(
    input dbus_req_t cache_dreq,
    output dbus_resp_t cache_dresp
);
    
endmodule